-------------------------------------------------------------------------------
-- Title      : Testbench for Fetch
-- Project    : 
-------------------------------------------------------------------------------
-- File       : Test_Fetch.vhd
-- Author     : Robert Jarzmik  <robert.jarzmik@free.fr>
-- Company    : 
-- Created    : 2016-11-11
-- Last update: 2016-11-11
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Testbench for Fetch
-------------------------------------------------------------------------------
-- Copyright (c) 2016 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2016-11-11  1.0      rj      Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity Test_Fetch is

  generic (
    );

  port (
    );

end entity Test_Fetch;

-------------------------------------------------------------------------------

architecture only of Test_Fetch is

  -----------------------------------------------------------------------------
  -- Internal signal declarations
  -----------------------------------------------------------------------------
  component Fetch
    port (
      
      );
  end component;

  signal clk   : bit := '0';
  signal reset : bit := '0';

begin  -- architecture str


  dut : Fetch port map (
    );
  -----------------------------------------------------------------------------
  -- Component instantiations
  -----------------------------------------------------------------------------

end architecture str;

-------------------------------------------------------------------------------

